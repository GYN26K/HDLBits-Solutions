module top_module(
    input clk,
    input load,
    input [255:0] data,
    output [255:0] q ); 

    wire [15:0] k [15:0] ; 

    

endmodule

// Alternate solution as systemVerilog has 2 D vectors availble where Verilog doesnt 