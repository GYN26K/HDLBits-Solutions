module top_module ( input a, input b, output out );
    
    mod_a an (a , b , out);

endmodule
