module top_module(
    input clk,
    input load,
    input [255:0] data,
    output [255:0] q ); 

endmodule