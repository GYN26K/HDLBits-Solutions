module top_module(
    input clk,
    input [7:0] in,
    input reset,    // Synchronous reset
    output done); //

    // State transition logic (combinational)

    // State flip-flops (sequential)
 
    // Output logic

endmodule 